module writeback();
endmodule
