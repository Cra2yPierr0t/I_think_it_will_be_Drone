module uart_top(
        input   logic RX,
        output  logic TX,
    );
    
endmodule
