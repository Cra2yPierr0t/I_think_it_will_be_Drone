module core_v0();

endmodule
